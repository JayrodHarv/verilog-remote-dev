`timescale 1ns/1ps

module beans (
    // input clk,
    // input rst
);

    // reg / wire declarations here

    // always @(posedge clk) begin
    // end

endmodule
