`timescale 1ns/1ps

module e (
    
);

    // reg / wire declarations here


endmodule
